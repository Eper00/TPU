module Floating_point_Unit#(
    parameter DATA_WIDTH = 16
)(
    input wire clk,                 
    input wire reset,                
    input wire en,
    input wire dec,    
    input wire [DATA_WIDTH-1:0] a,
    input wire [DATA_WIDTH-1:0] b,
    output reg [DATA_WIDTH-1:0] result
);

reg [4:0] a_exponent, b_exponent, result_exponent;
reg [9:0] a_fraction, b_fraction, result_fraction;
reg a_sign, b_sign, result_sign;
reg [21:0] product_fraction; // Szorzás után nagyobb méret kell
reg [5:0] shift_amount; // Maximum exponenskülönbség 31 lehet, ezért 6 bit elég
reg [11:0] extended_a_fraction, extended_b_fraction; // Mantissza + implicit 1 bit + extra hely shifteléshez
reg [11:0] sum_fraction;

always @(posedge clk or posedge reset) begin
    if (reset) begin
        result_exponent <= 0;
        result_fraction <= 0;
        result_sign <= 0;
        product_fraction<=0;
        shift_amount<=0; // Maximum exponenskülönbség 31 lehet, ezért 6 bit elég
        extended_a_fraction<=0; 
        extended_b_fraction<=0; // Mantissza + implicit 1 bit + extra hely shifteléshez
        sum_fraction<=0;
    end else if (en) begin
       

        if (dec == 0) begin
           // **ÖSSZEADÁS**
            

            if (a_exponent > b_exponent) begin
                result_exponent <= a_exponent;
                shift_amount = a_exponent - b_exponent;
                extended_b_fraction = {1'b1, b_fraction} >> shift_amount; // Jobbra shift a kisebb exponenshez
                extended_a_fraction = {1'b1, a_fraction}; // Nagyobb szám marad változatlanul
            end else begin
                result_exponent = b_exponent;
                shift_amount = b_exponent - a_exponent;
                extended_a_fraction = {1'b1, a_fraction} >> shift_amount; 
                extended_b_fraction = {1'b1, b_fraction}; 
            end

            // Mantisszák összeadása
            if (a_sign==b_sign)begin
                sum_fraction = extended_a_fraction + extended_b_fraction;
                if (a_sign==0)begin
                result_sign=0;
                end
                else begin
                result_sign=1;
                end
            end else begin
                if (a_sign==0)begin
                    if (extended_a_fraction>=extended_b_fraction)begin
                    sum_fraction = extended_a_fraction - extended_b_fraction;
                    result_sign=0;
                    end else begin 
                    sum_fraction = -1*extended_a_fraction + extended_b_fraction;
                    result_sign=1;
                    end
                    
                end else begin
                   if (extended_a_fraction>=extended_b_fraction)begin
                    sum_fraction = extended_a_fraction - extended_b_fraction;
                    result_sign=1;
                    end else begin 
                    sum_fraction = -1*extended_a_fraction + extended_b_fraction;
                    result_sign=0;
                    end
                    
                end
            end
            

            // **Normalizáció**
            if (sum_fraction[11]) begin
                result_fraction = sum_fraction[10:1]; // Ha túlcsordul, 1 bitet le kell shiftelni
                result_exponent = result_exponent + 1; // Kitevő növelése
            end else begin
                result_fraction = sum_fraction[9:0]; // Normál 10 bit
            end

            result_sign = a_sign; // Az előjel az erősebb számé marad

            
        end else begin
            // *** SZORZÁS ***
            result_sign = a_sign ^ b_sign;
            result_exponent = a_exponent + b_exponent - 15;
            product_fraction = {1,a_fraction} * {1,b_fraction};
           
            // Normalizálás
            if (product_fraction[21]) begin
                result_fraction = product_fraction[20:11];
                result_exponent = result_exponent + 1;
            end else begin
                result_fraction = product_fraction[19:10];
            end
             if (a==0||b==0)begin
                result_sign=0;
                result_exponent=0; 
                result_fraction=0;
            end
        end
    end
end
 // Bitek szétválasztása
  assign a_sign     = a[15];
  assign a_exponent = a[14:10];
  assign a_fraction = a[9:0]; // Implicit 1-es bit hozzáadása
  assign b_sign     = b[15];
  assign b_exponent = b[14:10];
  assign b_fraction = b[9:0]; // Implicit 1-es bit hozzáadása


assign result = {result_sign, result_exponent, result_fraction};

endmodule
